//Header file where we define a enum type for the instructions, ti identify better the
//executing instruction in the waveform of the modelsim.
enum {
    _add  ,
    _addu ,
    _and  ,
    _jr   ,
    _nor  ,
    _or   ,
    _slt  ,
    _sltu ,
    _sll  ,
    _srl  ,
    _sub  ,
    _subu ,
    _addi ,
    _addiu,
    _andi ,
    _beq  ,
    _bne  ,
    _lbu  ,
    _lhu  ,
    _ll   ,
    _lui  ,
    _lw   ,
    _ori  ,
    _slti ,
    _sltiu,
    _sb   ,
    _sc   ,
    _sh   ,
    _sw   ,
    _j    ,
    _jal  ,
    _mul  ,
    _nop
} INSTR;